* ADG1236 MACROMODEL
* Description: Converter
* Generic Desc: +/- 15V DUAL SPDT LOW CAP I.C.
* Developed by: Y.WONG 
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (09/2008)
* Copyright 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model 
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include: 
*
* END Notes
*
* Connections
*      1  = IN1
*      2  = S1A
*      3  = D1
*      4  = S1B 
*      5  = VSS
*      6  = GND
*      7  = NC
*      8  = NC
*      9  = IN2
*      10 = S2A
*      11 = D2
*      12 = S2B
*      13 = VDD
*      14 = NC
*      15 = NC
*      16 = NC
*****************
.SUBCKT ADG1236 1 2 3 4 5 6 9 10 11 12 13

X1 2 3 1 13 6 5 HIGHONSWITCH
X2 4 3 1 13 6 5 LOWONSWITCH
X3 10 11 9 13 6 5 HIGHONSWITCH
X4 12 11 9 13 6 5 LOWONSWITCH
DIN1A 1 13 DX
DIN1B 6 1 DX
DIN2A 9 13 DX
DIN2B 6 9 DX
CIN1 1 6 2p
CIN2 9 6 2p
CC1A1B 2 4 0.11p
CC2A2B 10 12 0.11p
CC1A2A 2 10 0.11p
CC1B2B 4 12 0.11p
RC1A2A 2 10 1.413E6
RC1B2B 4 12 1.413E6

.MODEL DX D(IS=1E-12 N=0.5 RS=0.1)
.ENDS

****************
* Logic Low On Switch
*
* Connections
*      101 = S
*      102 = D
*      103 = VIN
*      104 = VDD 
*      105 = GND
*      106 = VSS
*****************

.SUBCKT LOWONSWITCH  101 102 103 104 105 106

x1 103 104 105 107 NOTGATE
X2 107 108 104 106 105 VSENSE
X3 108 105 109 ENABLEDELAY
X4 101 102 109 104 105 106 SWITCH

*MODELS USED
.ENDS

****************
* Logic High On Switch
*
* Connections
*      101 = S
*      102 = D
*      103 = VIN
*      104 = VDD 
*      105 = GND
*      106 = VSS
*****************

.SUBCKT HIGHONSWITCH  101 102 103 104 105 106
x1 103 104 105 107 BUFF
X2 107 108 104 106 105 VSENSE
X3 108 105 109 ENABLEDELAY
X4 101 102 109 104 105 106 SWITCH

*MODELS USED
.ENDS

*****************
* NOT LOGIC
*
* Connections
*      201 = INPUT
*      202 = VDD
*      203 = GND
*      204 = OUTPUT
*****************
.SUBCKT NOTGATE 201 202 203 204

SNOT 205 203 201 203 SMOD2
RNOT 205 202 5G
EBUFFER 204 203 205 203 1

*MODELS USED
.MODEL SMOD2 VSWITCH(RON=1E-3 ROFF=1E11 VON=2.0 VOFF=0.8)
.ENDS


*****************
* BUFF LOGIC
*
* Connections
*      201 = INPUT
*      202 = VDD
*      203 = GND
*      204 = OUTPUT
*****************
.SUBCKT BUFF 201 202 203 204
SBUFF 205 203 201 203 SMOD2
RBUFF 205 202 5G
EBUFFER 204 203 205 203 1

*MODELS USED
.MODEL SMOD2 VSWITCH(RON=1E-3 ROFF=1E11 VON=0.8 VOFF=2.0)
.ENDS

****************
* Switch
*
* Connections
*      201 = S
*      202 = D
*      203 = VIN
*      204 = VDD 
*      205 = GND
*      206 = VSS
*****************

.SUBCKT SWITCH  201 202 203 204 205 206

*ANALOG SWITCH
S1 201 208 203 205 SMOD1
S2 204 207 203 205 SMOD2
S3 204 223 201 205 SMOD3 
S4 204 224 202 205 SMOD3
S5 223 207 201 205 SMOD7
S6 224 207 202 205 SMOD7
RD 207 205 5G
S7 208 202 207 205 SMOD4

DS1 201 204 DX 
DS2 206 201 DX
DD1 202 204 DX
DD2 206 202 DX

*ON OFF ISOLATION*
CSD 201 202 0.637p

*BANDWIDTH  
CSB 201 204 1.0p
CDB 202 204 1.0p

*CHARGE INJECTION
CGS 201 203 0.09p
CGD 202 203 0.09p

*MODELS USED
.MODEL SMOD1 VSWITCH(RON=120 ROFF=7.905E5 VON=2.0 VOFF=0.8)
.MODEL SMOD2 VSWITCH(RON=1E-3 ROFF=1E11 VON=2.0 VOFF=0.8)
.MODEL SMOD3 VSWITCH(RON=1E-3 ROFF=1E11 VON=0.8 VOFF=1.0)
.MODEL SMOD4 VSWITCH(RON=1E-3 ROFF=10E11 VON=4 VOFF=3)
.MODEL SMOD7 VSWITCH(RON=1E-3 ROFF=1E11 VON=-0.8 VOFF=-1.0)
.MODEL DX D(IS=1E-12 N=0.5 RS=0.1)
.ENDS

*****************
* ENABLE DELAY
*
* Connections
*      301 = INPUT
*      302 = COM
*      303 = OUTPUT
*****************
.SUBCKT ENABLEDELAY 301 302 303

EENBUFFER 304 302 301 302 1
RFEN 304 306 170k
CFEN 306 302 5p
DBREAKEN 306 305 DZ
RBEN 305 304 9k
EENBUFFEROUT 303 302 306 302 1 

*MODELS USED
.MODEL DZ D(IS=1E-14 N=0.04)
.ENDS

*****************
* OPERATING VOLTAGE 
*
* Connections
*      601 = INPUT
*      602 = OUTPUT
*      603 = VDD
*      604 = VSS
*      605 = GND
*****************
.SUBCKT VSENSE 601 602 603 604 605
SD1 601 606 603 605 SMOD3
SD2 606 607 603 605 SMOD4
SD3 607 608 605 604 SMOD5
SD4 608 609 605 604 SMOD6
RD0 609 605 5G
EBUFFER 602 605 609 605 1

*MODELS USED
.MODEL SMOD3 VSWITCH(RON=1E-3 ROFF=1E11 VON=12.0 VOFF=11.9)
.MODEL SMOD4 VSWITCH(RON=1E-3 ROFF=1E11 VON=16.5 VOFF=16.6)
.MODEL SMOD5 VSWITCH(RON=1E-3 ROFF=1E11 VON=0 VOFF=-0.1)
.MODEL SMOD6 VSWITCH(RON=1E-3 ROFF=1E11 VON=16.5 VOFF=16.6)
.ENDS







