* ADG659 MACROMODEL MODEL CAN ONLY RUN ON SPICE2
* Description: Converter
* Generic Desc: 3V/5V  4/8 Channel Analog muxs
* Developed by: Y.WONG 
* Revision History: 08/10/2012 - Updated to new header style
* 1.1 (11/2008)
* Copyright 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model 
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include: 
*
* END Notes
*
* Connections
*      1  = S1B
*      2  = S3B
*      3  = DB
*      4  = S4B 
*      5  = S2B
*      6  = /EN
*      7  = VSS
*      8  = GND
*      9  = A1
*      10 = A0
*      11 = S4A
*      12 = S1A
*      13 = DA
*      14 = S2A
*      15 = S3A
*      16 = VDD
*****************
.SUBCKT ADG659 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
RL1 16 8 5000MEG
RL2 7 8 5000MEG
CEN 6 8 2p
CA0 10 8 2p
CA1 9 8 2p
DENA 6 16 DY
DENB 7 6 DY
DA0A 10 16 DY
DA0B 7 10 DY
DA1A 9 16 DY
DA1B 7 9 DY
X9 6 10 9 16 8 17 18 19 20 DECODER
X1 12 13 17 16 8 7 6 HIGHONSWITCH
X2 14 13 18 16 8 7 6 HIGHONSWITCH
X3 15 13 19 16 8 7 6 HIGHONSWITCH
X4 11 13 20 16 8 7 6  HIGHONSWITCH
X5 1 3 17 16 8 7 6  HIGHONSWITCH
X6 5 3 18 16 8 7 6  HIGHONSWITCH
X7 2 3 19 16 8 7 6  HIGHONSWITCH
X8 4 3 20 16 8 7 6  HIGHONSWITCH
CS12 12 14 0.15p
CS13 12 15 0.15p
CS14 12 11 0.15p
CS15 12 1 0.15p
CS16 12 5 0.15p
CS17 12 2 0.15p
CS18 12 4 0.15p
CS23 14 15 0.15p
CS24 14 11 0.15p
CS25 14 1 0.15p
CS26 14 5 0.15p
CS27 14 2 0.15p
CS28 14 4 0.15p
CS34 15 11 0.15p
CS35 15 1 0.15p
CS36 15 5 0.15p
CS37 15 2 0.15p
CS38 15 4 0.15p
CS45 11 1 0.15p
CS46 11 5 0.15p
CS47 11 2 0.15p
CS48 11 4 0.15p
CS56 1 5 0.15p
CS57 1 2 0.15p
CS58 1 4 0.15p
CS67 5 2 0.15p
CS68 5 4 0.15p
CS78 2 4 0.15p
*MODELS USED
.MODEL DY D(IS=1E-14 N=0.04 RS=30)
.ENDS
*****************
* 2 to 4 with Enable Decoder
*
* Connections
*      101 = /EN
*      102 = A0
*      103 = A1
*      104 = VDD 
*      105 = GND
*      106 = D1
*      107 = D2
*      108 = D3
*      109 = D4
*****************

.SUBCKT DECODER 101 102 103 104 105 106 107 108 109
SEN 124 105 101 105 SMOD2
SA0 110 105 102 105 SMOD2
SA1 111 105 103 105 SMOD2
SD1A 104 112 124 105 SMOD2
SD1B 112 113 110 105 SMOD2
SD1C 113 114 111 105 SMOD2
SD2A 104 115 124 105 SMOD2
SD2B 115 116 102 105 SMOD2
SD2C 116 117 111 105 SMOD2
SD3A 104 118 124 105 SMOD2
SD3B 118 119 110 105 SMOD2
SD3C 119 120 103 105 SMOD2
SD4A 104 121 124 105 SMOD2
SD4B 121 122 102 105 SMOD2
SD4C 122 123 103 105 SMOD2
REN 124 104 5G
RA0 110 104 5G
RA1 111 104 5G
RD1 105 114 5G
RD2 105 117 5G
RD3 105 120 5G
RD4 105 123 5G
ED1 106 105 114 105 1
ED2 107 105 117 105 1
ED3 108 105 120 105 1
ED4 109 105 123 105 1

*MODELS USED
.MODEL SMOD2 VSWITCH(RON=1E-3 ROFF=1E11 VON=2.0 VOFF=0.8)
.ENDS

****************
* Logic High On Switch
*
* Connections
*      101 = S
*      102 = D
*      103 = VIN
*      104 = VDD 
*      105 = GND
*      106 = VSS
*      107 = /EN
*****************

.SUBCKT HIGHONSWITCH  101 102 103 104 105 106 107

x1 103 104 105 108 BUFF
X2 108 109 104 106 105 VSENSE
X3 109 110 107 105 ENABLE
X4 110 105 111 ENABLEDELAY
X5 101 102 111 104 105 106 SWITCH

*MODELS USED
.ENDS

****************
* Switch
*
* Connections
*      201 = S
*      202 = D
*      203 = VIN
*      204 = VDD 
*      205 = GND
*      206 = VSS
*****************

.SUBCKT SWITCH  201 202 203 204 205 206

*ANALOG SWITCH
EBuffer 214 205 202 205 1
S1 210 202 203 205 SMOD1
Vo2 214 219 0
EVDD 219 220 204 205 1
SN 210 209 205 220 SMOD7
Vo1 205 218 0
EVSS 217 218 206 205 1
SP 210 208 214 217 SMOD8 
Xn 215 209 214 205 204 206 VCRN
Xp 207 208 214 205 204 206 VCRP
RS1 201 207 1
RS2 201 215 1

DS1 201 204 DX 
DS2 206 201 DX
DD1 202 204 DX
DD2 206 202 DX

*ON OFF ISOLATION*
CSD 201 202 0.201p
 
*BANDWIDTH * 
CSB 201 206 2.1p
CDB 202 204 2.1p

*CHARGE INJECTION
CGS 201 203 0.167p
CGD 202 203 0.167p

*MODELS USED
.MODEL SMOD1 VSWITCH(RON=1 ROFF=7E11 VON=2.0 VOFF=0.8)
.MODEL SMOD7 VSWITCH(RON=1E-3 ROFF=1E11 VON=0.81 VOFF=0.79)
.MODEL SMOD8 VSWITCH(RON=1E-3 ROFF=1E11 VON=1.21 VOFF=1.19)
.MODEL DX D(IS=1E-12 N=0.04 RS=120)
.ENDS

*****************
* BUFF LOGIC
*
* Connections
*      201 = INPUT
*      202 = VDD
*      203 = GND
*      204 = OUTPUT
*****************
.SUBCKT BUFF 201 202 203 204
SBUFF 205 203 201 203 SMOD2
RBUFF 205 202 5G
EBUFFER 204 203 205 203 1

*MODELS USED
.MODEL SMOD2 VSWITCH(RON=1E-3 ROFF=1E11 VON=0.8 VOFF=2.0)
.ENDS

*****************
* ENABLE DELAY
*
* Connections
*      301 = INPUT
*      302 = COM
*      303 = OUTPUT
*****************
.SUBCKT ENABLEDELAY 301 302 303

EENBUFFER 304 302 301 302 1
RFEN 304 306 45k
CFEN 306 302 5p
DBREAKEN 306 305 DZ
RBEN 305 304 17k
EENBUFFEROUT 303 302 306 302 1 

*MODELS USED
.MODEL DZ D(IS=1E-14 N=0.04)
.ENDS

*****************
* Enable ON/OFF 
*
* Connections
*      501 = INPUT
*      502 = OUTPUT
*      503 = VIN
*      504 = GND
*****************
.SUBCKT ENABLE 501 502 503 504 
SENABLE 501 505 503 504 SMOD2
RD0 505 504 5G
EBUFFER 502 504 505 504 1

*MODELS USED
.MODEL SMOD2 VSWITCH(RON=1E-3 ROFF=1E11 VON=0.8 VOFF=2.0)
.ENDS

*****************
* OPERATING VOLTAGE 
*
* Connections
*      601 = INPUT
*      602 = OUTPUT
*      603 = VDD
*      604 = VSS
*      605 = GND
*****************
.SUBCKT VSENSE 601 602 603 604 605
SD1 601 606 603 605 SMOD3
SD2 606 607 603 605 SMOD4
SD3 607 608 605 604 SMOD5
SD4 608 609 605 604 SMOD6
SD5 609 602 603 604 SMOD7
RD0 602 605 5G

*MODELS USED
.MODEL SMOD3 VSWITCH(RON=1E-3 ROFF=1E11 VON=2 VOFF=1.9)
.MODEL SMOD4 VSWITCH(RON=1E-3 ROFF=1E11 VON=12 VOFF=12.1)
.MODEL SMOD5 VSWITCH(RON=1E-3 ROFF=1E11 VON=0 VOFF=-0.1)
.MODEL SMOD6 VSWITCH(RON=1E-3 ROFF=1E11 VON=6 VOFF=6.1)
.MODEL SMOD7 VSWITCH(RON=1E-3 ROFF=1E11 VON=12 VOFF=12.1)

.ENDS

*****************
* Voltage Controlled Resistance n-channel
*
* Connections
*      701 = R+
*      702 = R-
*      704 = V+
*      705 = V-
*      707 = VDD
*      711 = VSS
*****************
.SUBCKT VCRN 701 702 704 705 707 711
vtn 708 0 0.8
ERES 701 703 VALUE={285*V(706,0)*(1/(V(707,0)-V(704,705)-V(708,0)))}
VSENSE 703 702 0
FCOPY 0 706 VSENSE 1
RRES 706 0 1
.ENDS

*****************
* Voltage Controlled Resistance p-channel
*
* Connections
*      701 = R+
*      702 = R-
*      704 = V+
*      705 = V-
*      707 = VDD
*      711 = VSS
*****************
.SUBCKT VCRP 701 702 704 705 707 711
vtp 708 0 1.2
ERES 701 703 VALUE={246*V(706,0)*(1/(V(704,705)-V(711,0)-V(708,0)))}
VSENSE 703 702 0
FCOPY 0 706 VSENSE 1
RRES 706 0 1
.ENDS




