* D:\Neuro repos\memristive-brain\test-circuits\LTSPICE\NON-memristor_neuron\multivibrator+\NE555 multivibrator+.asc
XU1 0 N002 N004 N001 N005 N002 N003 N001 NE555
C1 N001 0 100�F V=25
C2 N002 0 0.68�F V=25
R3 0 N006 10k tol=5
R2 N003 N002 4.3k tol=5
V1 N001 0 5
C3 N005 0 0.1�F
R1 N001 N003 5.1k tol=5
D2 N003 N002 1N4148
R4 N004 N006 10k tol=5
.model D D
.lib C:\Users\Alexe\Documents\LTspiceXVII\lib\cmp\standard.dio
.lib NE555.sub
.backanno
.end

