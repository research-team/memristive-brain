* ADG609 MACROMODEL
* Description: Converter
* Generic Desc: 3V dual 4-channel multiplexer
* Developed by: Y.WONG 
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (03/2008)
* Copyright 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model 
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include: 
*
* END Notes
*
* Connections
*      1  = A0
*      2  = EN
*      3  = VSS
*      4  = S1A 
*      5  = S2A
*      6  = S3A
*      7  = S4A
*      8  = DA
*      9  = DB
*      10 = S4B
*      11 = S3B
*      12 = S2B
*      13 = S1B
*      14 = VDD
*      15 = GND
*      16 = A1
*****************
.SUBCKT ADG609 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
RL1 14 15 100MEG
RL2 3 15 500MEG
DA0A 1 14 DY
DA0B 15 1 DY
DA1A 16 14 DY
DA1B 15 16 DY
DENA 2 14 DY
DENB 15 2 DY
CA0 1 15 5p
CA1 16 15 5p
CEN 2 15 5p
X5 2 17 14 3 15 VSENSE
X4 17 15 18 ENABLEDELAY
X2 1 15 19 ADDRESSDELAY
X3 16 15 20 ADDRESSDELAY
X1 18 19 20 14 15 21 22 23 24 DECODER
X6 21 15 25 BBMDELAY
X7 22 15 26 BBMDELAY
X8 23 15 27 BBMDELAY
X9 24 15 28 BBMDELAY
X10 4 8 25 14 15 3 SWITCH
X11 13 9 25 14 15 3 SWITCH
X12 5 8 26 14 15 3 SWITCH
X13 12 9 26 14 15 3 SWITCH
X14 6 8 27 14 15 3 SWITCH
X15 11 9 27 14 15 3 SWITCH
X21 7 8 28 14 15 3 SWITCH
X22 10 9 28 14 15 3 SWITCH
CS12A 4 5 0.01p
CS12B 13 12 0.01p
CS13A 4 6 0.01p
CS13B 13 11 0.01p
CS14A 4 7 0.01p
CS14B 13 10 0.01p
CS23A 5 6 0.01p
CS23B 12 11 0.01p
CS24A 5 7 0.01p
CS24B 12 10 0.01p
CS34A 6 7 0.01p
CS34B 11 10 0.01p

*MODELS USED
.MODEL DY D(IS=1E-14 N=0.04 RS=15)
.ENDS

*****************
* 2 to 4 with Enable Decoder
*
* Connections
*      101 = EN
*      102 = A0
*      103 = A1
*      104 = VDD 
*      105 = GND
*      106 = D1
*      107 = D2
*      108 = D3
*      109 = D4
*****************

.SUBCKT DECODER 101 102 103 104 105 106 107 108 109
SA0 110 105 102 105 SMOD2
SA1 111 105 103 105 SMOD2
SD1A 104 112 101 105 SMOD2
SD1B 112 113 110 105 SMOD2
SD1C 113 114 111 105 SMOD2
SD2A 104 115 101 105 SMOD2
SD2B 115 116 102 105 SMOD2
SD2C 116 117 111 105 SMOD2
SD3A 104 118 101 105 SMOD2
SD3B 118 119 110 105 SMOD2
SD3C 119 120 103 105 SMOD2
SD4A 104 121 101 105 SMOD2
SD4B 121 122 102 105 SMOD2
SD4C 122 123 103 105 SMOD2
RA0 110 104 33G
RA1 111 104 33G
RD1 105 114 33G
RD2 105 117 33G
RD3 105 120 33G
RD4 105 123 33G
ED1 106 105 114 105 1
ED2 107 105 117 105 1
ED3 108 105 120 105 1
ED4 109 105 123 105 1

*MODELS USED
.MODEL SMOD2 VSWITCH(RON=1E-3 ROFF=1E13 VON=2.4 VOFF=0.8)
.ENDS

****************
* Switch
*
* Connections
*      201 = S
*      202 = D
*      203 = VIN
*      204 = VDD 
*      205 = GND
*      206 = VSS
*****************

.SUBCKT SWITCH  201 202 203 204 205 206

*ANALOG SWITCH
S1 201 202 203 205 SMOD1

*LEAKAGE CuRRENT 
S2 201 207 202 201 SMOD2
S3 202 208 202 201 SMOD2
S4 201 209 202 201 SMOD3
S5 202 210 202 201 SMOD3
I1 207 205 8.61n
I2 205 208 8.61n
I3 205 209 8.61n
I4 210 205 8.61n

DS1 201 204 DX 
DS2 206 201 DX
DD1 202 204 DX
DD2 206 202 DX


*ON OFF ISOLATION*
CSD 201 202 0.087p

*BANDWIDTH * No Bandwidth Data
CSB 201 206 8.9p
CDB 202 204 4.9p

*CHARGE INJECTION
CGS 201 203 0.1p
CGD 202 203 0.1p

*MODELS USED
.MODEL SMOD1 VSWITCH(RON=40 ROFF=562E6 VON=2.4 VOFF=0.8)
.MODEL SMOD2 VSWITCH(RON=1E-03 ROFF=1E13 VON=2.2 VOFF=1.1)
.MODEL SMOD3 VSWITCH(RON=1E-03 ROFF=1E13 VON=-2.2 VOFF=-1.1)
.MODEL DX D(IS=1E-14 N=0.04 RS=15)
.ENDS

*****************
* ENABLE DELAY
*
* Connections
*      301 = INPUT
*      302 = COM
*      303 = OUTPUT
*****************
.SUBCKT ENABLEDELAY 301 302 303

EENBUFFER 304 302 301 302 1
RFEN 304 303 31k
CFEN 303 302 5p
DBREAKEN 303 305 DZ
RBEN 305 304 12.5k

*MODELS USED
.MODEL DZ D(IS=1E-14 N=0.04)
.ENDS

*****************
* ADDRESS DELAY
*
* Connections
*      401 = INPUT
*      402 = COM
*      403 = OUTPUT
*****************
.SUBCKT ADDRESSDELAY 401 402 403

EADBUFFER 404 402 401 402 1
RFAD 404 403 15k
CFAD 403 402 5p

*MODELS USED
.MODEL DZ D(IS=1E-14 N=1)
.ENDS

*****************
* BBM DELAY
*
* Connections
*      501 = INPUT
*      502 = COM
*      503 = OUTPUT
*****************
.SUBCKT BBMDELAY 501 502 503

RFBBM 501 504 3.2k
CFBBM 504 502 5p
DBREAKBBM 504 505 DZ
RBBBM 505 501 0
EBBMBUFFER 503 502 504 502 1

*MODELS USED
.MODEL DZ D(IS=1E-14 N=0.04)
.ENDS

*****************
* OPERATING VOLTAGE 
*
* Connections
*      601 = INPUT
*      602 = OUTPUT
*      603 = VDD
*      604 = VSS
*      605 = GND
*****************
.SUBCKT VSENSE 601 602 603 604 605
SD1 601 606 603 605 SMOD3
SD2 606 607 603 605 SMOD4
SD3 607 608 605 604 SMOD5
SD4 608 602 605 604 SMOD6
RD0 602 605 33G

*MODELS USED
.MODEL SMOD3 VSWITCH(RON=1E-3 ROFF=1E20 VON=2.7 VOFF=2.6)
.MODEL SMOD4 VSWITCH(RON=1E-3 ROFF=1E20 VON=5.5 VOFF=5.6)
.MODEL SMOD5 VSWITCH(RON=1E-3 ROFF=1E20 VON=0 VOFF=-0.1)
.MODEL SMOD6 VSWITCH(RON=1E-3 ROFF=1E20 VON=5.5 VOFF=5.6)

.ENDS



